
// gate level circuit
module and_2_gatelevel(output wire F,  input wire A, input wire B);
    and(F, A, B);
endmodule


//data_flow model
module and_2_data_flow(output wire F,  input wire A, input wire B);
    assign F = A & B;
endmodule


// Behavioural Model of the AND gate.
module and_2_behave(output reg F,  input wire A, input wire B);
    always @ (A or B) begin
        if ((A == 1'b1)  &  (B == 1'b1))
        begin
            F = 1'b1;
        end
        else
            F = 1'b0;
    end
endmodule  

module tb;
    reg A1,B1;
    wire F1;


    //and_2_gatelevel instance0(F1, A1, B1);
    //and_2_behave instance1(F1, A1, B1);
    and_2_data_flow instance2(F1, A1, B1);

    initial begin
        A1 = 0; B1 = 0;
        #1  A1 = 0; B1 = 1;
        #1  A1 = 1; B1 = 0;
        #1  A1 = 1; B1 = 1;
        #1;
    end

    initial begin
        $monitor("%t A1=%d, B1=%d, F1=%d" , $time, A1,B1,F1);
        $dumpfile("dump.vcd");
        $dumpvars();
    end
endmodule