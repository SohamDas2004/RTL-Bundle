// NOT Gate Modelling

// gate level circuit
module not_gatelevel(output wire F,  input wire A);
    not(F, A);
endmodule

//data_flow model
module not_data_flow(output wire F,  input wire A);
    assign F = ~A;
endmodule

// Behavioural Model of the AND gate.
module not_behave(output reg F,  input wire A);
    always @ (A ) begin
        if (A == 1'b0)
        begin
            F = 1'b1;
        end
        else
        begin
            F = 1'b0;
        end
    end
endmodule  

module tb;
    reg A0,A1,A2;
    wire F0,F1,F2;

    not_gatelevel instance0(F0, A0);
    not_data_flow instance1(F1, A1);
    not_behave instance2(F2, A2);

    initial begin
        A0 = 0;A1=1;A2=0;
        #1  A0 = 1;A1=0;A2=1;
        #1;
    end

    initial begin
        $display("NOT  gate circuit");
        $monitor("%t A0=%d,F0=%d , A1=%d,F1=%d, A2=%d,F2=%d" ,$time, A0,F0,A1,F1,A2,F2);
        $dumpfile("dump.vcd");
        $dumpvars();
    end
endmodule